
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity subtractor is
    port (
    );
end subtractor;

architecture arch of subtractor is

begin


end arch;
